import_C("tEV3Platform.h");

celltype tEV3Platform{
	entry sTaskBody eTaskBody;
};
